module XORR (input logic sinal_1, sinal_2, output logic Xor_out);	
		assign Xor_out = sinal_1 ^ sinal_2;	
endmodule: XORR